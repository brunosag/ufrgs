library verilog;
use verilog.vl_types.all;
entity rca4_vlg_vec_tst is
end rca4_vlg_vec_tst;
