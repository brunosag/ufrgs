library verilog;
use verilog.vl_types.all;
entity fa_vlg_vec_tst is
end fa_vlg_vec_tst;
