library verilog;
use verilog.vl_types.all;
entity rca_vlg_vec_tst is
end rca_vlg_vec_tst;
